module ram_controller(); 